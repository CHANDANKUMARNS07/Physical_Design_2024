VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO avsdpll
  CLASS BLOCK ;
  FOREIGN avsdpll ;
  ORIGIN 0.000 0.000 ;
  SIZE 36.180 BY 13.710 ;
  SITE unithddb1 ;
  PIN GND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 10.030 10.380 10.250 10.970 ;
        RECT 11.590 10.380 11.760 11.170 ;
        RECT 14.250 10.380 14.420 11.160 ;
        RECT 16.980 10.380 17.150 11.170 ;
        RECT 18.090 10.380 18.260 11.170 ;
        RECT 9.320 10.210 18.670 10.380 ;
        RECT 0.990 9.740 10.340 9.910 ;
        RECT 11.400 9.740 20.750 9.910 ;
        RECT 1.700 9.150 1.920 9.740 ;
        RECT 3.260 8.950 3.430 9.740 ;
        RECT 5.920 8.960 6.090 9.740 ;
        RECT 8.650 8.950 8.820 9.740 ;
        RECT 9.760 8.950 9.930 9.740 ;
        RECT 12.110 9.150 12.330 9.740 ;
        RECT 13.670 8.950 13.840 9.740 ;
        RECT 16.330 8.960 16.500 9.740 ;
        RECT 19.060 8.950 19.230 9.740 ;
        RECT 20.170 8.950 20.340 9.740 ;
      LAYER mcon ;
        RECT 9.670 10.210 9.840 10.380 ;
        RECT 10.510 10.210 10.680 10.380 ;
        RECT 11.350 10.210 11.520 10.380 ;
        RECT 12.530 10.210 12.700 10.380 ;
        RECT 13.370 10.210 13.540 10.380 ;
        RECT 14.430 10.210 14.600 10.380 ;
        RECT 15.350 10.210 15.520 10.380 ;
        RECT 16.700 10.210 16.870 10.380 ;
        RECT 17.500 10.210 17.670 10.380 ;
        RECT 18.340 10.210 18.510 10.380 ;
        RECT 1.340 9.740 1.510 9.910 ;
        RECT 2.180 9.740 2.350 9.910 ;
        RECT 3.020 9.740 3.190 9.910 ;
        RECT 4.200 9.740 4.370 9.910 ;
        RECT 5.040 9.740 5.210 9.910 ;
        RECT 6.100 9.740 6.270 9.910 ;
        RECT 7.020 9.740 7.190 9.910 ;
        RECT 8.370 9.740 8.540 9.910 ;
        RECT 9.170 9.740 9.340 9.910 ;
        RECT 10.010 9.740 10.180 9.910 ;
        RECT 11.750 9.740 11.920 9.910 ;
        RECT 12.590 9.740 12.760 9.910 ;
        RECT 13.430 9.740 13.600 9.910 ;
        RECT 14.610 9.740 14.780 9.910 ;
        RECT 15.450 9.740 15.620 9.910 ;
        RECT 16.510 9.740 16.680 9.910 ;
        RECT 17.430 9.740 17.600 9.910 ;
        RECT 18.780 9.740 18.950 9.910 ;
        RECT 19.580 9.740 19.750 9.910 ;
        RECT 20.420 9.740 20.590 9.910 ;
      LAYER met1 ;
        RECT 9.320 10.060 18.670 10.540 ;
        RECT 0.000 9.750 0.310 9.890 ;
        RECT 0.590 9.750 10.340 10.060 ;
        RECT 0.000 9.580 10.340 9.750 ;
        RECT 11.400 9.580 20.750 10.060 ;
        RECT 0.000 9.120 0.900 9.580 ;
        RECT 0.000 8.980 0.310 9.120 ;
    END
  END GND
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 21.140 9.820 34.410 10.910 ;
        RECT 2.480 8.510 3.550 8.580 ;
        RECT 2.480 8.460 3.670 8.510 ;
        RECT 1.020 8.220 3.670 8.460 ;
        RECT 5.240 8.220 6.380 8.570 ;
        RECT 1.020 8.210 6.380 8.220 ;
        RECT 7.970 8.560 11.450 8.570 ;
        RECT 12.890 8.560 13.960 8.580 ;
        RECT 21.140 8.570 26.420 9.820 ;
        RECT 29.420 9.810 34.410 9.820 ;
        RECT 30.710 8.760 34.410 9.810 ;
        RECT 31.070 8.750 34.410 8.760 ;
        RECT 7.970 8.510 13.960 8.560 ;
        RECT 7.970 8.220 14.080 8.510 ;
        RECT 15.650 8.220 16.790 8.570 ;
        RECT 7.970 8.210 16.790 8.220 ;
        RECT 18.380 8.210 26.420 8.570 ;
        RECT 1.020 6.860 26.420 8.210 ;
        RECT 1.900 6.720 26.420 6.860 ;
        RECT 1.900 5.810 29.330 6.720 ;
        RECT 2.380 5.250 29.330 5.810 ;
        RECT 6.060 5.130 29.330 5.250 ;
        RECT 6.060 5.060 16.830 5.130 ;
        RECT 8.790 4.820 16.830 5.060 ;
        RECT 10.630 4.690 16.830 4.820 ;
        RECT 10.970 4.540 16.830 4.690 ;
        RECT 11.080 4.490 16.830 4.540 ;
        RECT 20.250 4.390 29.330 5.130 ;
        RECT 20.250 4.350 28.090 4.390 ;
        RECT 20.250 4.340 21.550 4.350 ;
        RECT 20.250 4.040 21.180 4.340 ;
      LAYER li1 ;
        RECT 33.940 8.930 34.110 10.240 ;
        RECT 1.700 7.230 1.930 7.840 ;
        RECT 3.260 7.230 3.430 8.330 ;
        RECT 5.920 7.230 6.090 8.340 ;
        RECT 8.650 7.230 8.820 8.330 ;
        RECT 9.760 7.230 9.930 8.330 ;
        RECT 12.110 7.230 12.340 7.840 ;
        RECT 13.670 7.230 13.840 8.330 ;
        RECT 16.330 7.230 16.500 8.340 ;
        RECT 19.060 7.230 19.230 8.330 ;
        RECT 20.170 7.230 20.340 8.330 ;
        RECT 1.020 7.040 10.340 7.230 ;
        RECT 11.430 7.040 20.750 7.230 ;
        RECT 23.360 7.210 23.700 7.990 ;
        RECT 21.140 7.040 30.160 7.210 ;
        RECT 8.470 6.680 29.330 6.700 ;
        RECT 1.010 6.530 29.330 6.680 ;
        RECT 1.010 6.510 8.680 6.530 ;
        RECT 2.660 6.180 3.080 6.510 ;
        RECT 2.520 5.970 3.230 6.180 ;
        RECT 6.780 5.540 7.010 6.510 ;
        RECT 11.150 6.310 29.150 6.530 ;
        RECT 22.050 4.660 28.820 4.870 ;
      LAYER mcon ;
        RECT 1.610 7.040 1.800 7.230 ;
        RECT 2.470 7.040 2.660 7.230 ;
        RECT 3.330 7.040 3.520 7.230 ;
        RECT 4.530 7.040 4.720 7.230 ;
        RECT 5.610 7.040 5.800 7.230 ;
        RECT 6.550 7.040 6.740 7.230 ;
        RECT 7.330 7.040 7.520 7.230 ;
        RECT 8.780 7.040 8.970 7.230 ;
        RECT 9.600 7.040 9.790 7.230 ;
        RECT 12.020 7.040 12.210 7.230 ;
        RECT 12.880 7.040 13.070 7.230 ;
        RECT 13.740 7.040 13.930 7.230 ;
        RECT 14.940 7.040 15.130 7.230 ;
        RECT 16.020 7.040 16.210 7.230 ;
        RECT 16.960 7.040 17.150 7.230 ;
        RECT 17.740 7.040 17.930 7.230 ;
        RECT 19.190 7.040 19.380 7.230 ;
        RECT 20.010 7.040 20.200 7.230 ;
        RECT 21.370 7.040 21.540 7.210 ;
        RECT 21.710 7.040 21.880 7.210 ;
        RECT 22.050 7.040 22.220 7.210 ;
        RECT 22.390 7.040 22.560 7.210 ;
        RECT 22.730 7.040 22.900 7.210 ;
        RECT 23.070 7.040 23.240 7.210 ;
        RECT 23.410 7.040 23.580 7.210 ;
        RECT 23.750 7.040 23.920 7.210 ;
        RECT 24.090 7.040 24.260 7.210 ;
        RECT 24.430 7.040 24.600 7.210 ;
        RECT 24.770 7.040 24.940 7.210 ;
        RECT 25.110 7.040 25.280 7.210 ;
        RECT 25.450 7.040 25.620 7.210 ;
        RECT 25.790 7.040 25.960 7.210 ;
        RECT 26.130 7.040 26.300 7.210 ;
        RECT 26.470 7.040 26.640 7.210 ;
        RECT 26.810 7.040 26.980 7.210 ;
        RECT 27.150 7.040 27.320 7.210 ;
        RECT 27.490 7.040 27.660 7.210 ;
        RECT 27.830 7.040 28.000 7.210 ;
        RECT 28.170 7.040 28.340 7.210 ;
        RECT 28.510 7.040 28.680 7.210 ;
        RECT 28.850 7.040 29.020 7.210 ;
        RECT 29.190 7.040 29.360 7.210 ;
        RECT 29.530 7.040 29.700 7.210 ;
        RECT 29.870 7.040 30.040 7.210 ;
        RECT 1.810 6.510 1.980 6.680 ;
        RECT 2.150 6.510 2.320 6.680 ;
        RECT 2.490 6.510 2.660 6.680 ;
        RECT 2.830 6.510 3.000 6.680 ;
        RECT 3.170 6.510 3.340 6.680 ;
        RECT 3.510 6.510 3.680 6.680 ;
        RECT 3.850 6.510 4.020 6.680 ;
        RECT 4.190 6.510 4.360 6.680 ;
        RECT 4.530 6.510 4.700 6.680 ;
        RECT 4.870 6.510 5.040 6.680 ;
        RECT 5.210 6.510 5.380 6.680 ;
        RECT 5.550 6.510 5.720 6.680 ;
        RECT 5.890 6.510 6.060 6.680 ;
        RECT 6.230 6.510 6.400 6.680 ;
        RECT 6.570 6.510 6.740 6.680 ;
        RECT 6.910 6.510 7.080 6.680 ;
        RECT 7.250 6.510 7.420 6.680 ;
        RECT 7.590 6.510 7.760 6.680 ;
        RECT 8.880 6.530 9.050 6.700 ;
        RECT 9.220 6.530 9.390 6.700 ;
        RECT 9.560 6.530 9.730 6.700 ;
        RECT 9.900 6.530 10.070 6.700 ;
        RECT 10.240 6.530 10.410 6.700 ;
        RECT 10.580 6.530 10.750 6.700 ;
        RECT 10.920 6.530 11.090 6.700 ;
        RECT 11.260 6.530 11.430 6.700 ;
        RECT 11.600 6.530 11.770 6.700 ;
        RECT 11.940 6.530 12.110 6.700 ;
        RECT 12.280 6.530 12.450 6.700 ;
        RECT 12.620 6.530 12.790 6.700 ;
        RECT 12.960 6.530 13.130 6.700 ;
        RECT 13.300 6.530 13.470 6.700 ;
        RECT 13.640 6.530 13.810 6.700 ;
        RECT 13.980 6.530 14.150 6.700 ;
        RECT 14.320 6.530 14.490 6.700 ;
        RECT 14.660 6.530 14.830 6.700 ;
        RECT 15.000 6.530 15.170 6.700 ;
        RECT 15.340 6.530 15.510 6.700 ;
        RECT 15.680 6.530 15.850 6.700 ;
        RECT 16.020 6.530 16.190 6.700 ;
        RECT 16.360 6.530 16.530 6.700 ;
        RECT 16.700 6.530 16.870 6.700 ;
        RECT 17.040 6.530 17.210 6.700 ;
        RECT 17.380 6.530 17.550 6.700 ;
        RECT 17.720 6.530 17.890 6.700 ;
        RECT 18.060 6.530 18.230 6.700 ;
        RECT 18.400 6.530 18.570 6.700 ;
        RECT 18.740 6.530 18.910 6.700 ;
        RECT 19.080 6.530 19.250 6.700 ;
        RECT 19.420 6.530 19.590 6.700 ;
        RECT 19.760 6.530 19.930 6.700 ;
        RECT 20.100 6.530 20.270 6.700 ;
        RECT 20.440 6.530 20.610 6.700 ;
        RECT 20.780 6.530 20.950 6.700 ;
        RECT 21.120 6.530 21.290 6.700 ;
        RECT 21.460 6.530 21.630 6.700 ;
        RECT 21.800 6.530 21.970 6.700 ;
        RECT 22.140 6.530 22.310 6.700 ;
        RECT 22.480 6.530 22.650 6.700 ;
        RECT 22.820 6.530 22.990 6.700 ;
        RECT 23.160 6.530 23.330 6.700 ;
        RECT 23.500 6.530 23.670 6.700 ;
        RECT 23.840 6.530 24.010 6.700 ;
        RECT 24.180 6.530 24.350 6.700 ;
        RECT 24.520 6.530 24.690 6.700 ;
        RECT 24.860 6.530 25.030 6.700 ;
        RECT 25.200 6.530 25.370 6.700 ;
        RECT 25.540 6.530 25.710 6.700 ;
        RECT 25.880 6.530 26.050 6.700 ;
        RECT 26.220 6.530 26.390 6.700 ;
        RECT 26.560 6.530 26.730 6.700 ;
        RECT 26.900 6.530 27.070 6.700 ;
        RECT 27.240 6.530 27.410 6.700 ;
        RECT 27.580 6.530 27.750 6.700 ;
        RECT 27.920 6.530 28.090 6.700 ;
        RECT 28.260 6.530 28.430 6.700 ;
        RECT 28.600 6.530 28.770 6.700 ;
        RECT 28.940 6.530 29.110 6.700 ;
        RECT 27.490 4.680 27.660 4.850 ;
        RECT 27.920 4.680 28.090 4.850 ;
      LAYER met1 ;
        RECT 0.000 7.340 0.310 7.410 ;
        RECT 0.000 6.860 10.340 7.340 ;
        RECT 11.430 7.030 20.750 7.340 ;
        RECT 21.140 7.030 30.160 7.340 ;
        RECT 11.430 6.860 30.160 7.030 ;
        RECT 0.000 6.670 29.330 6.860 ;
        RECT 0.000 6.500 0.320 6.670 ;
        RECT 1.010 6.380 29.330 6.670 ;
        RECT 27.430 4.920 28.130 6.380 ;
        RECT 27.430 4.620 28.150 4.920 ;
    END
  END VDD
  PIN ENb_CP
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 3.024000 ;
    PORT
      LAYER li1 ;
        RECT 31.440 9.940 31.770 10.110 ;
        RECT 32.570 7.660 32.900 7.870 ;
        RECT 33.440 7.680 33.770 7.850 ;
        RECT 8.740 5.520 9.100 5.610 ;
        RECT 8.740 5.510 9.610 5.520 ;
        RECT 8.740 5.270 9.630 5.510 ;
        RECT 8.740 5.260 9.610 5.270 ;
        RECT 8.740 5.250 9.100 5.260 ;
      LAYER mcon ;
        RECT 31.520 9.940 31.690 10.110 ;
        RECT 32.650 7.680 32.820 7.850 ;
        RECT 33.520 7.680 33.690 7.850 ;
        RECT 8.770 5.340 8.940 5.510 ;
      LAYER met1 ;
        RECT 31.450 9.860 31.770 10.180 ;
        RECT 32.580 7.910 32.900 7.920 ;
        RECT 32.580 7.610 34.530 7.910 ;
        RECT 32.580 7.600 32.900 7.610 ;
        RECT 8.690 5.250 9.040 5.610 ;
      LAYER via ;
        RECT 31.480 9.890 31.740 10.150 ;
        RECT 32.610 7.630 32.870 7.890 ;
        RECT 8.720 5.280 9.010 5.570 ;
      LAYER met2 ;
        RECT 31.450 10.140 31.770 10.180 ;
        RECT 31.450 9.890 32.300 10.140 ;
        RECT 31.450 9.860 31.770 9.890 ;
        RECT 32.050 8.940 32.300 9.890 ;
        RECT 31.820 8.700 32.300 8.940 ;
        RECT 32.050 7.910 32.300 8.700 ;
        RECT 32.580 7.910 32.900 7.920 ;
        RECT 32.050 7.610 32.900 7.910 ;
        RECT 32.580 7.600 32.900 7.610 ;
        RECT 32.590 7.450 32.870 7.600 ;
        RECT 28.720 7.150 32.890 7.450 ;
        RECT 28.720 7.030 29.250 7.150 ;
        RECT 3.020 6.710 29.250 7.030 ;
        RECT 0.000 5.840 0.280 6.060 ;
        RECT 3.020 5.840 3.350 6.710 ;
        RECT 0.000 5.520 3.350 5.840 ;
        RECT 0.000 5.290 0.280 5.520 ;
        RECT 8.690 5.250 9.040 6.710 ;
    END
  END ENb_CP
  PIN CLK
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.351000 ;
    ANTENNADIFFAREA 0.469800 ;
    PORT
      LAYER li1 ;
        RECT 12.010 12.220 12.180 12.560 ;
        RECT 20.300 11.770 20.680 11.850 ;
        RECT 20.300 11.540 20.690 11.770 ;
        RECT 18.010 11.370 20.760 11.540 ;
        RECT 20.210 11.180 20.760 11.370 ;
        RECT 21.380 11.180 21.550 11.930 ;
        RECT 15.970 10.800 16.300 10.980 ;
        RECT 20.210 10.950 21.550 11.180 ;
        RECT 20.210 10.940 21.210 10.950 ;
        RECT 21.380 9.650 21.550 10.950 ;
      LAYER mcon ;
        RECT 12.010 12.300 12.180 12.470 ;
        RECT 20.420 11.570 20.590 11.740 ;
        RECT 18.090 11.370 18.260 11.540 ;
        RECT 16.050 10.810 16.220 10.980 ;
      LAYER met1 ;
        RECT 11.950 12.550 12.230 12.560 ;
        RECT 11.950 12.130 12.240 12.550 ;
        RECT 17.100 12.240 18.320 12.560 ;
        RECT 17.100 12.130 17.350 12.240 ;
        RECT 11.950 11.880 17.350 12.130 ;
        RECT 18.030 11.330 18.320 12.240 ;
        RECT 20.340 11.500 20.660 11.820 ;
        RECT 18.030 11.040 18.310 11.330 ;
        RECT 15.960 10.750 18.310 11.040 ;
      LAYER via ;
        RECT 20.370 11.530 20.630 11.790 ;
      LAYER met2 ;
        RECT 20.310 11.470 20.690 11.850 ;
        RECT 29.190 1.570 29.920 1.920 ;
        RECT 29.190 1.140 30.340 1.570 ;
        RECT 29.810 0.280 30.340 1.140 ;
        RECT 29.690 0.000 30.460 0.280 ;
      LAYER via2 ;
        RECT 20.360 11.520 20.640 11.800 ;
        RECT 29.250 1.200 29.850 1.860 ;
      LAYER met3 ;
        RECT 20.310 11.570 20.930 11.850 ;
        RECT 20.310 11.470 20.940 11.570 ;
        RECT 20.550 5.550 20.940 11.470 ;
        RECT 20.550 5.540 22.930 5.550 ;
        RECT 20.550 5.140 23.300 5.540 ;
        RECT 22.680 4.370 23.300 5.140 ;
        RECT 22.680 2.300 23.310 4.370 ;
        RECT 22.690 1.610 23.310 2.300 ;
        RECT 29.190 1.610 29.920 1.920 ;
        RECT 22.690 1.130 29.920 1.610 ;
    END
  END CLK
  PIN ENb_VCO
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.063000 ;
    PORT
      LAYER li1 ;
        RECT 23.350 8.360 23.700 8.700 ;
      LAYER mcon ;
        RECT 23.440 8.460 23.610 8.630 ;
      LAYER met1 ;
        RECT 21.260 8.380 23.670 8.690 ;
        RECT 21.360 8.100 21.800 8.380 ;
      LAYER via ;
        RECT 21.410 8.150 21.670 8.410 ;
      LAYER met2 ;
        RECT 2.890 10.200 19.740 10.210 ;
        RECT 2.890 9.920 21.720 10.200 ;
        RECT 0.000 8.280 0.280 8.540 ;
        RECT 2.890 8.280 3.200 9.920 ;
        RECT 18.040 9.910 21.720 9.920 ;
        RECT 21.380 8.460 21.720 9.910 ;
        RECT 0.000 7.990 3.200 8.280 ;
        RECT 21.360 8.090 21.720 8.460 ;
        RECT 0.000 7.770 0.280 7.990 ;
    END
  END ENb_VCO
  PIN GND#2
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 5.350 3.750 6.020 4.560 ;
        RECT 6.790 3.820 7.010 4.340 ;
        RECT 6.570 3.750 7.240 3.820 ;
        RECT 5.350 3.730 8.850 3.750 ;
        RECT 9.970 3.730 15.040 4.010 ;
        RECT 17.270 3.730 17.690 3.980 ;
        RECT 5.350 3.580 19.080 3.730 ;
        RECT 8.680 3.560 19.080 3.580 ;
        RECT 19.810 3.560 29.330 3.730 ;
        RECT 1.790 3.220 2.000 3.240 ;
        RECT 1.710 3.050 2.070 3.220 ;
        RECT 1.790 2.970 2.000 3.050 ;
        RECT 9.600 2.500 9.790 3.560 ;
        RECT 10.840 2.500 11.030 3.560 ;
        RECT 12.680 3.190 17.920 3.560 ;
        RECT 20.750 3.280 28.240 3.560 ;
        RECT 12.680 3.180 18.090 3.190 ;
        RECT 12.550 3.010 18.090 3.180 ;
        RECT 13.290 3.000 18.090 3.010 ;
        RECT 2.740 1.380 2.920 1.740 ;
        RECT 7.040 1.160 7.260 1.490 ;
      LAYER mcon ;
        RECT 5.950 3.580 6.120 3.750 ;
        RECT 6.290 3.580 6.460 3.750 ;
        RECT 6.630 3.580 6.800 3.750 ;
        RECT 6.970 3.580 7.140 3.750 ;
        RECT 7.310 3.580 7.480 3.750 ;
        RECT 7.650 3.580 7.820 3.750 ;
        RECT 8.880 3.560 9.050 3.730 ;
        RECT 9.220 3.560 9.390 3.730 ;
        RECT 9.560 3.560 9.730 3.730 ;
        RECT 9.900 3.560 10.070 3.730 ;
        RECT 10.240 3.560 10.410 3.730 ;
        RECT 10.580 3.560 10.750 3.730 ;
        RECT 10.920 3.560 11.090 3.730 ;
        RECT 11.260 3.560 11.430 3.730 ;
        RECT 11.600 3.560 11.770 3.730 ;
        RECT 11.940 3.560 12.110 3.730 ;
        RECT 12.280 3.560 12.450 3.730 ;
        RECT 12.620 3.560 12.790 3.730 ;
        RECT 12.960 3.560 13.130 3.730 ;
        RECT 13.300 3.560 13.470 3.730 ;
        RECT 13.640 3.560 13.810 3.730 ;
        RECT 13.980 3.560 14.150 3.730 ;
        RECT 14.320 3.560 14.490 3.730 ;
        RECT 14.660 3.560 14.830 3.730 ;
        RECT 15.000 3.560 15.170 3.730 ;
        RECT 15.340 3.560 15.510 3.730 ;
        RECT 15.680 3.560 15.850 3.730 ;
        RECT 16.020 3.560 16.190 3.730 ;
        RECT 16.360 3.560 16.530 3.730 ;
        RECT 16.700 3.560 16.870 3.730 ;
        RECT 17.040 3.560 17.210 3.730 ;
        RECT 17.380 3.560 17.550 3.730 ;
        RECT 17.720 3.560 17.890 3.730 ;
        RECT 18.060 3.560 18.230 3.730 ;
        RECT 18.400 3.560 18.570 3.730 ;
        RECT 18.740 3.560 18.910 3.730 ;
        RECT 20.100 3.560 20.270 3.730 ;
        RECT 20.440 3.560 20.610 3.730 ;
        RECT 20.780 3.560 20.950 3.730 ;
        RECT 21.120 3.560 21.290 3.730 ;
        RECT 21.460 3.560 21.630 3.730 ;
        RECT 21.800 3.560 21.970 3.730 ;
        RECT 22.140 3.560 22.310 3.730 ;
        RECT 22.480 3.560 22.650 3.730 ;
        RECT 22.820 3.560 22.990 3.730 ;
        RECT 23.160 3.560 23.330 3.730 ;
        RECT 23.500 3.560 23.670 3.730 ;
        RECT 23.840 3.560 24.010 3.730 ;
        RECT 24.180 3.560 24.350 3.730 ;
        RECT 24.520 3.560 24.690 3.730 ;
        RECT 24.860 3.560 25.030 3.730 ;
        RECT 25.200 3.560 25.370 3.730 ;
        RECT 25.540 3.560 25.710 3.730 ;
        RECT 25.880 3.560 26.050 3.730 ;
        RECT 26.220 3.560 26.390 3.730 ;
        RECT 26.560 3.560 26.730 3.730 ;
        RECT 26.900 3.560 27.070 3.730 ;
        RECT 27.240 3.560 27.410 3.730 ;
        RECT 27.580 3.560 27.750 3.730 ;
        RECT 27.920 3.560 28.090 3.730 ;
        RECT 28.260 3.560 28.430 3.730 ;
        RECT 28.600 3.560 28.770 3.730 ;
        RECT 1.810 3.050 1.980 3.220 ;
        RECT 2.750 1.470 2.920 1.640 ;
        RECT 7.080 1.240 7.250 1.410 ;
      LAYER met1 ;
        RECT 0.000 4.660 0.310 4.830 ;
        RECT 0.000 4.230 1.020 4.660 ;
        RECT 0.000 3.920 0.310 4.230 ;
        RECT 0.650 3.900 1.020 4.230 ;
        RECT 0.650 3.420 29.330 3.900 ;
        RECT 1.750 2.990 2.050 3.420 ;
        RECT 3.290 1.700 3.530 3.420 ;
        RECT 2.690 1.410 3.530 1.700 ;
        RECT 6.610 1.470 6.880 3.420 ;
        RECT 6.610 1.180 7.280 1.470 ;
    END
  END GND#2
  PIN VDD#2
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 7.780 3.530 8.930 3.540 ;
        RECT 5.440 3.410 8.930 3.530 ;
        RECT 4.980 2.140 8.930 3.410 ;
        RECT 4.980 2.030 11.820 2.140 ;
        RECT 4.980 0.770 6.150 2.030 ;
        RECT 8.090 1.630 11.820 2.030 ;
        RECT 8.090 0.780 12.570 1.630 ;
        RECT 19.220 1.610 20.060 2.060 ;
        RECT 19.220 0.770 21.080 1.610 ;
      LAYER li1 ;
        RECT 7.030 3.000 7.260 3.390 ;
        RECT 8.050 3.120 8.460 3.290 ;
        RECT 7.030 2.710 7.340 3.000 ;
        RECT 8.110 2.830 8.410 3.120 ;
        RECT 7.030 2.690 7.260 2.710 ;
        RECT 8.050 2.660 8.460 2.830 ;
        RECT 8.110 2.390 8.410 2.660 ;
        RECT 8.050 2.220 8.460 2.390 ;
        RECT 5.700 0.770 5.910 1.880 ;
        RECT 11.890 0.780 12.570 1.190 ;
        RECT 20.270 0.780 21.080 1.280 ;
        RECT 8.470 0.770 29.340 0.780 ;
        RECT 1.010 0.610 29.340 0.770 ;
        RECT 1.010 0.600 8.680 0.610 ;
      LAYER mcon ;
        RECT 7.170 2.770 7.340 2.940 ;
        RECT 8.150 2.640 8.360 2.850 ;
        RECT 1.810 0.600 1.980 0.770 ;
        RECT 2.150 0.600 2.320 0.770 ;
        RECT 2.490 0.600 2.660 0.770 ;
        RECT 2.830 0.600 3.000 0.770 ;
        RECT 3.170 0.600 3.340 0.770 ;
        RECT 3.510 0.600 3.680 0.770 ;
        RECT 3.850 0.600 4.020 0.770 ;
        RECT 4.190 0.600 4.360 0.770 ;
        RECT 4.530 0.600 4.700 0.770 ;
        RECT 4.870 0.600 5.040 0.770 ;
        RECT 5.210 0.600 5.380 0.770 ;
        RECT 5.550 0.600 5.720 0.770 ;
        RECT 5.890 0.600 6.060 0.770 ;
        RECT 6.230 0.600 6.400 0.770 ;
        RECT 6.570 0.600 6.740 0.770 ;
        RECT 6.910 0.600 7.080 0.770 ;
        RECT 7.250 0.600 7.420 0.770 ;
        RECT 7.590 0.600 7.760 0.770 ;
        RECT 8.880 0.610 9.050 0.780 ;
        RECT 9.220 0.610 9.390 0.780 ;
        RECT 9.560 0.610 9.730 0.780 ;
        RECT 9.900 0.610 10.070 0.780 ;
        RECT 10.240 0.610 10.410 0.780 ;
        RECT 10.580 0.610 10.750 0.780 ;
        RECT 10.920 0.610 11.090 0.780 ;
        RECT 11.260 0.610 11.430 0.780 ;
        RECT 11.600 0.610 11.770 0.780 ;
        RECT 11.940 0.610 12.110 0.780 ;
        RECT 12.280 0.610 12.450 0.780 ;
        RECT 12.620 0.610 12.790 0.780 ;
        RECT 12.960 0.610 13.130 0.780 ;
        RECT 13.300 0.610 13.470 0.780 ;
        RECT 13.640 0.610 13.810 0.780 ;
        RECT 13.980 0.610 14.150 0.780 ;
        RECT 14.320 0.610 14.490 0.780 ;
        RECT 14.660 0.610 14.830 0.780 ;
        RECT 15.000 0.610 15.170 0.780 ;
        RECT 15.340 0.610 15.510 0.780 ;
        RECT 15.680 0.610 15.850 0.780 ;
        RECT 16.020 0.610 16.190 0.780 ;
        RECT 16.360 0.610 16.530 0.780 ;
        RECT 16.700 0.610 16.870 0.780 ;
        RECT 17.040 0.610 17.210 0.780 ;
        RECT 17.380 0.610 17.550 0.780 ;
        RECT 17.720 0.610 17.890 0.780 ;
        RECT 18.060 0.610 18.230 0.780 ;
        RECT 18.400 0.610 18.570 0.780 ;
        RECT 18.740 0.610 18.910 0.780 ;
        RECT 19.080 0.610 19.250 0.780 ;
        RECT 19.420 0.610 19.590 0.780 ;
        RECT 19.760 0.610 19.930 0.780 ;
        RECT 20.100 0.610 20.270 0.780 ;
        RECT 20.440 0.610 20.610 0.780 ;
        RECT 20.780 0.610 20.950 0.780 ;
        RECT 21.120 0.610 21.290 0.780 ;
        RECT 21.460 0.610 21.630 0.780 ;
        RECT 21.800 0.610 21.970 0.780 ;
        RECT 22.140 0.610 22.310 0.780 ;
        RECT 22.480 0.610 22.650 0.780 ;
        RECT 22.820 0.610 22.990 0.780 ;
        RECT 23.160 0.610 23.330 0.780 ;
        RECT 23.500 0.610 23.670 0.780 ;
        RECT 23.840 0.610 24.010 0.780 ;
        RECT 24.180 0.610 24.350 0.780 ;
        RECT 24.520 0.610 24.690 0.780 ;
        RECT 24.860 0.610 25.030 0.780 ;
        RECT 25.200 0.610 25.370 0.780 ;
        RECT 25.540 0.610 25.710 0.780 ;
        RECT 25.880 0.610 26.050 0.780 ;
        RECT 26.220 0.610 26.390 0.780 ;
        RECT 26.560 0.610 26.730 0.780 ;
        RECT 26.900 0.610 27.070 0.780 ;
        RECT 27.240 0.610 27.410 0.780 ;
        RECT 27.580 0.610 27.750 0.780 ;
        RECT 27.920 0.610 28.090 0.780 ;
        RECT 28.260 0.610 28.430 0.780 ;
        RECT 28.600 0.610 28.770 0.780 ;
      LAYER met1 ;
        RECT 7.110 2.710 8.420 3.000 ;
        RECT 7.570 2.530 8.420 2.710 ;
        RECT 7.570 0.940 7.870 2.530 ;
        RECT 1.010 0.460 29.340 0.940 ;
        RECT 28.530 0.310 29.040 0.460 ;
        RECT 28.320 0.000 29.230 0.310 ;
    END
  END VDD#2
  PIN VCO_IN
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.313200 ;
    PORT
      LAYER li1 ;
        RECT 32.880 8.800 33.050 9.650 ;
        RECT 32.880 8.530 33.200 8.800 ;
        RECT 32.880 8.050 33.050 8.530 ;
      LAYER mcon ;
        RECT 33.010 8.570 33.180 8.740 ;
      LAYER met1 ;
        RECT 35.210 8.810 35.530 8.820 ;
        RECT 32.950 8.510 35.530 8.810 ;
        RECT 35.210 8.500 35.530 8.510 ;
      LAYER via ;
        RECT 35.240 8.530 35.500 8.790 ;
      LAYER met2 ;
        RECT 35.900 8.820 36.180 9.040 ;
        RECT 35.210 8.500 36.180 8.820 ;
        RECT 35.900 8.270 36.180 8.500 ;
    END
  END VCO_IN
  PIN VDD#3
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER nwell ;
        RECT 9.350 11.910 18.670 13.260 ;
        RECT 9.350 11.900 14.710 11.910 ;
        RECT 9.350 11.660 12.000 11.900 ;
        RECT 10.810 11.610 12.000 11.660 ;
        RECT 10.810 11.540 11.880 11.610 ;
        RECT 13.570 11.550 14.710 11.900 ;
        RECT 16.300 11.550 18.670 11.910 ;
      LAYER li1 ;
        RECT 9.350 12.890 18.670 13.080 ;
        RECT 20.180 12.940 30.160 13.110 ;
        RECT 10.030 12.280 10.260 12.890 ;
        RECT 11.590 11.790 11.760 12.890 ;
        RECT 14.250 11.780 14.420 12.890 ;
        RECT 16.980 11.790 17.150 12.890 ;
        RECT 18.090 11.790 18.260 12.890 ;
      LAYER mcon ;
        RECT 9.940 12.890 10.130 13.080 ;
        RECT 10.800 12.890 10.990 13.080 ;
        RECT 11.660 12.890 11.850 13.080 ;
        RECT 12.860 12.890 13.050 13.080 ;
        RECT 13.940 12.890 14.130 13.080 ;
        RECT 14.880 12.890 15.070 13.080 ;
        RECT 15.660 12.890 15.850 13.080 ;
        RECT 17.110 12.890 17.300 13.080 ;
        RECT 17.930 12.890 18.120 13.080 ;
        RECT 20.350 12.940 20.520 13.110 ;
        RECT 20.690 12.940 20.860 13.110 ;
        RECT 21.030 12.940 21.200 13.110 ;
        RECT 21.370 12.940 21.540 13.110 ;
        RECT 21.710 12.940 21.880 13.110 ;
        RECT 22.050 12.940 22.220 13.110 ;
        RECT 22.390 12.940 22.560 13.110 ;
        RECT 22.730 12.940 22.900 13.110 ;
        RECT 23.070 12.940 23.240 13.110 ;
        RECT 23.410 12.940 23.580 13.110 ;
        RECT 23.750 12.940 23.920 13.110 ;
        RECT 24.090 12.940 24.260 13.110 ;
        RECT 24.430 12.940 24.600 13.110 ;
        RECT 24.770 12.940 24.940 13.110 ;
        RECT 25.110 12.940 25.280 13.110 ;
        RECT 25.450 12.940 25.620 13.110 ;
        RECT 25.790 12.940 25.960 13.110 ;
        RECT 26.130 12.940 26.300 13.110 ;
        RECT 26.470 12.940 26.640 13.110 ;
        RECT 26.810 12.940 26.980 13.110 ;
        RECT 27.150 12.940 27.320 13.110 ;
        RECT 27.490 12.940 27.660 13.110 ;
        RECT 27.830 12.940 28.000 13.110 ;
        RECT 28.170 12.940 28.340 13.110 ;
        RECT 28.510 12.940 28.680 13.110 ;
        RECT 28.850 12.940 29.020 13.110 ;
        RECT 29.190 12.940 29.360 13.110 ;
        RECT 29.530 12.940 29.700 13.110 ;
        RECT 29.870 12.940 30.040 13.110 ;
      LAYER met1 ;
        RECT 18.420 13.260 21.630 13.270 ;
        RECT 9.350 12.780 32.170 13.260 ;
        RECT 31.380 11.650 32.170 12.780 ;
        RECT 31.380 11.640 35.600 11.650 ;
        RECT 31.380 11.240 35.620 11.640 ;
        RECT 31.380 11.230 35.130 11.240 ;
        RECT 35.280 9.960 35.620 11.240 ;
        RECT 35.870 9.960 36.180 10.180 ;
        RECT 35.280 9.340 36.180 9.960 ;
        RECT 35.870 9.270 36.180 9.340 ;
    END
  END VDD#3
  PIN REF
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.879000 ;
    ANTENNADIFFAREA 0.214500 ;
    PORT
      LAYER li1 ;
        RECT 3.430 5.980 4.530 6.170 ;
        RECT 3.430 5.670 3.660 5.980 ;
        RECT 1.050 2.200 1.320 3.970 ;
        RECT 1.050 1.910 3.110 2.200 ;
        RECT 1.570 1.570 1.950 1.910 ;
      LAYER mcon ;
        RECT 1.680 1.670 1.850 1.840 ;
      LAYER met1 ;
        RECT 1.600 1.600 1.920 1.920 ;
      LAYER via ;
        RECT 1.630 1.630 1.890 1.890 ;
      LAYER met2 ;
        RECT 19.180 13.430 19.950 13.710 ;
        RECT 19.420 12.780 19.700 13.430 ;
        RECT 19.370 12.410 19.750 12.780 ;
        RECT 1.570 1.570 1.950 1.950 ;
      LAYER via2 ;
        RECT 19.420 12.450 19.700 12.730 ;
        RECT 1.620 1.620 1.900 1.900 ;
      LAYER met3 ;
        RECT 7.250 12.440 19.790 12.820 ;
        RECT 7.250 10.970 7.630 12.440 ;
        RECT 19.340 12.360 19.790 12.440 ;
        RECT 7.250 9.980 7.640 10.970 ;
        RECT 5.010 9.870 7.640 9.980 ;
        RECT 5.010 9.600 7.630 9.870 ;
        RECT 5.010 4.350 5.390 9.600 ;
        RECT 3.370 3.970 5.390 4.350 ;
        RECT 3.370 1.950 3.750 3.970 ;
        RECT 1.570 1.570 3.750 1.950 ;
    END
  END REF
  OBS
      LAYER li1 ;
        RECT 9.580 12.610 9.760 12.650 ;
        RECT 9.470 11.870 9.760 12.610 ;
        RECT 10.550 12.070 10.770 12.650 ;
        RECT 9.930 11.900 10.770 12.070 ;
        RECT 9.470 11.700 9.720 11.870 ;
        RECT 9.930 11.700 10.120 11.900 ;
        RECT 9.280 11.310 9.650 11.700 ;
        RECT 9.900 11.410 10.120 11.700 ;
        RECT 10.320 11.480 10.660 11.650 ;
        RECT 11.150 11.620 11.320 12.510 ;
        RECT 12.470 11.940 12.640 12.510 ;
        RECT 9.900 11.360 10.130 11.410 ;
        RECT 9.950 11.310 10.130 11.360 ;
        RECT 10.980 11.320 11.320 11.620 ;
        RECT 12.100 11.690 12.640 11.940 ;
        RECT 11.550 11.580 11.880 11.590 ;
        RECT 12.100 11.580 12.290 11.690 ;
        RECT 11.550 11.540 12.290 11.580 ;
        RECT 11.510 11.370 12.290 11.540 ;
        RECT 11.550 11.340 12.290 11.370 ;
        RECT 9.470 11.040 9.640 11.310 ;
        RECT 9.950 11.140 10.780 11.310 ;
        RECT 9.470 10.680 9.770 11.040 ;
        RECT 10.560 10.680 10.780 11.140 ;
        RECT 11.150 10.810 11.320 11.320 ;
        RECT 12.100 11.070 12.290 11.340 ;
        RECT 12.010 10.760 12.290 11.070 ;
        RECT 12.470 10.880 12.640 11.690 ;
        RECT 12.910 11.970 13.080 12.510 ;
        RECT 12.910 11.680 13.580 11.970 ;
        RECT 12.910 10.880 13.080 11.680 ;
        RECT 13.300 11.620 13.580 11.680 ;
        RECT 13.810 11.620 13.980 12.500 ;
        RECT 15.120 11.960 15.290 12.520 ;
        RECT 13.300 11.330 13.980 11.620 ;
        RECT 14.590 11.690 15.290 11.960 ;
        RECT 14.590 11.600 14.760 11.690 ;
        RECT 14.550 11.580 14.760 11.600 ;
        RECT 14.210 11.530 14.760 11.580 ;
        RECT 14.170 11.360 14.760 11.530 ;
        RECT 14.210 11.330 14.760 11.360 ;
        RECT 13.250 10.770 13.580 10.940 ;
        RECT 13.810 10.800 13.980 11.330 ;
        RECT 15.120 10.890 15.290 11.690 ;
        RECT 15.560 11.990 15.730 12.520 ;
        RECT 16.060 12.280 16.230 12.610 ;
        RECT 15.560 11.690 16.280 11.990 ;
        RECT 15.560 10.890 15.730 11.690 ;
        RECT 16.030 11.630 16.280 11.690 ;
        RECT 16.540 11.630 16.710 12.510 ;
        RECT 16.030 11.330 16.710 11.630 ;
        RECT 17.650 11.620 17.820 12.510 ;
        RECT 16.900 11.370 17.240 11.540 ;
        RECT 16.540 10.810 16.710 11.330 ;
        RECT 17.520 11.320 17.820 11.620 ;
        RECT 21.820 11.390 21.990 11.930 ;
        RECT 17.650 10.810 17.820 11.320 ;
        RECT 22.400 11.210 22.570 12.490 ;
        RECT 22.840 12.360 23.010 12.490 ;
        RECT 22.840 12.310 23.160 12.360 ;
        RECT 22.840 11.990 29.950 12.310 ;
        RECT 22.840 11.930 23.160 11.990 ;
        RECT 22.840 11.400 23.010 11.930 ;
        RECT 21.730 10.920 22.570 11.210 ;
        RECT 23.400 11.150 23.570 11.820 ;
        RECT 23.840 11.400 24.010 11.990 ;
        RECT 24.400 11.150 24.570 11.820 ;
        RECT 24.840 11.400 25.010 11.990 ;
        RECT 25.400 11.150 25.570 11.820 ;
        RECT 25.840 11.400 26.010 11.990 ;
        RECT 26.400 11.150 26.570 11.820 ;
        RECT 26.840 11.400 27.010 11.990 ;
        RECT 27.400 11.150 27.570 11.820 ;
        RECT 27.840 11.400 28.010 11.990 ;
        RECT 28.400 11.150 28.570 11.820 ;
        RECT 28.840 11.400 29.010 11.990 ;
        RECT 22.740 10.980 23.570 11.150 ;
        RECT 23.740 10.980 24.570 11.150 ;
        RECT 24.740 10.980 25.570 11.150 ;
        RECT 25.740 10.980 26.570 11.150 ;
        RECT 26.740 10.980 27.570 11.150 ;
        RECT 27.740 10.980 28.570 11.150 ;
        RECT 28.740 10.980 29.340 11.150 ;
        RECT 19.440 10.550 19.790 10.840 ;
        RECT 19.440 10.380 21.140 10.550 ;
        RECT 1.140 9.080 1.440 9.440 ;
        RECT 1.140 8.800 1.310 9.080 ;
        RECT 2.230 8.980 2.450 9.440 ;
        RECT 0.540 8.520 1.310 8.800 ;
        RECT 1.620 8.810 2.450 8.980 ;
        RECT 1.620 8.760 1.800 8.810 ;
        RECT 2.820 8.800 2.990 9.310 ;
        RECT 3.680 9.050 3.960 9.360 ;
        RECT 0.540 2.750 0.820 8.520 ;
        RECT 1.140 8.420 1.310 8.520 ;
        RECT 1.570 8.710 1.800 8.760 ;
        RECT 1.570 8.420 1.790 8.710 ;
        RECT 1.990 8.470 2.330 8.640 ;
        RECT 2.650 8.500 2.990 8.800 ;
        RECT 3.770 8.780 3.960 9.050 ;
        RECT 3.220 8.750 3.960 8.780 ;
        RECT 3.180 8.580 3.960 8.750 ;
        RECT 3.220 8.540 3.960 8.580 ;
        RECT 3.220 8.530 3.550 8.540 ;
        RECT 1.140 8.250 1.390 8.420 ;
        RECT 1.140 7.510 1.430 8.250 ;
        RECT 1.600 8.220 1.790 8.420 ;
        RECT 1.600 8.050 2.440 8.220 ;
        RECT 1.250 7.470 1.430 7.510 ;
        RECT 2.220 7.470 2.440 8.050 ;
        RECT 2.820 7.610 2.990 8.500 ;
        RECT 3.770 8.430 3.960 8.540 ;
        RECT 4.140 8.430 4.310 9.240 ;
        RECT 3.770 8.180 4.310 8.430 ;
        RECT 3.680 7.560 3.850 7.900 ;
        RECT 4.140 7.610 4.310 8.180 ;
        RECT 4.580 8.440 4.750 9.240 ;
        RECT 4.920 9.180 5.250 9.350 ;
        RECT 5.480 8.790 5.650 9.320 ;
        RECT 4.970 8.500 5.650 8.790 ;
        RECT 5.880 8.760 6.430 8.790 ;
        RECT 5.840 8.590 6.430 8.760 ;
        RECT 5.880 8.540 6.430 8.590 ;
        RECT 6.220 8.520 6.430 8.540 ;
        RECT 4.970 8.440 5.250 8.500 ;
        RECT 4.580 8.150 5.250 8.440 ;
        RECT 4.580 7.610 4.750 8.150 ;
        RECT 5.480 7.620 5.650 8.500 ;
        RECT 6.260 8.430 6.430 8.520 ;
        RECT 6.790 8.430 6.960 9.230 ;
        RECT 6.260 8.160 6.960 8.430 ;
        RECT 6.790 7.600 6.960 8.160 ;
        RECT 7.230 8.430 7.400 9.230 ;
        RECT 7.640 9.140 7.970 9.320 ;
        RECT 8.210 8.790 8.380 9.310 ;
        RECT 9.320 8.800 9.490 9.310 ;
        RECT 7.700 8.490 8.380 8.790 ;
        RECT 8.570 8.580 8.910 8.750 ;
        RECT 9.190 8.500 9.490 8.800 ;
        RECT 11.550 9.080 11.850 9.440 ;
        RECT 9.680 8.580 10.560 8.750 ;
        RECT 7.700 8.430 7.950 8.490 ;
        RECT 7.230 8.130 7.950 8.430 ;
        RECT 7.230 7.600 7.400 8.130 ;
        RECT 7.730 7.510 7.900 7.840 ;
        RECT 8.210 7.610 8.380 8.490 ;
        RECT 9.320 7.610 9.490 8.500 ;
        RECT 10.230 8.340 10.560 8.580 ;
        RECT 11.550 8.420 11.720 9.080 ;
        RECT 12.640 8.980 12.860 9.440 ;
        RECT 12.030 8.810 12.860 8.980 ;
        RECT 12.030 8.760 12.210 8.810 ;
        RECT 13.230 8.800 13.400 9.310 ;
        RECT 14.090 9.050 14.370 9.360 ;
        RECT 11.980 8.710 12.210 8.760 ;
        RECT 11.980 8.420 12.200 8.710 ;
        RECT 12.400 8.470 12.740 8.640 ;
        RECT 13.060 8.500 13.400 8.800 ;
        RECT 14.180 8.780 14.370 9.050 ;
        RECT 13.630 8.750 14.370 8.780 ;
        RECT 13.590 8.580 14.370 8.750 ;
        RECT 13.630 8.540 14.370 8.580 ;
        RECT 13.630 8.530 13.960 8.540 ;
        RECT 11.550 8.340 11.800 8.420 ;
        RECT 10.230 8.250 11.800 8.340 ;
        RECT 10.230 8.170 11.840 8.250 ;
        RECT 11.550 7.510 11.840 8.170 ;
        RECT 12.010 8.220 12.200 8.420 ;
        RECT 12.010 8.050 12.850 8.220 ;
        RECT 11.660 7.470 11.840 7.510 ;
        RECT 12.630 7.470 12.850 8.050 ;
        RECT 13.230 7.610 13.400 8.500 ;
        RECT 14.180 8.430 14.370 8.540 ;
        RECT 14.550 8.430 14.720 9.240 ;
        RECT 14.180 8.180 14.720 8.430 ;
        RECT 14.090 7.560 14.260 7.900 ;
        RECT 14.550 7.610 14.720 8.180 ;
        RECT 14.990 8.440 15.160 9.240 ;
        RECT 15.330 9.180 15.660 9.350 ;
        RECT 15.890 8.790 16.060 9.320 ;
        RECT 15.380 8.500 16.060 8.790 ;
        RECT 16.290 8.760 16.840 8.790 ;
        RECT 16.250 8.590 16.840 8.760 ;
        RECT 16.290 8.540 16.840 8.590 ;
        RECT 16.630 8.520 16.840 8.540 ;
        RECT 15.380 8.440 15.660 8.500 ;
        RECT 14.990 8.150 15.660 8.440 ;
        RECT 14.990 7.610 15.160 8.150 ;
        RECT 15.890 7.620 16.060 8.500 ;
        RECT 16.670 8.430 16.840 8.520 ;
        RECT 17.200 8.430 17.370 9.230 ;
        RECT 16.670 8.160 17.370 8.430 ;
        RECT 17.200 7.600 17.370 8.160 ;
        RECT 17.640 8.430 17.810 9.230 ;
        RECT 18.050 9.140 18.380 9.320 ;
        RECT 18.620 8.790 18.790 9.310 ;
        RECT 19.730 8.800 19.900 9.310 ;
        RECT 18.110 8.490 18.790 8.790 ;
        RECT 18.980 8.580 19.320 8.750 ;
        RECT 19.600 8.500 19.900 8.800 ;
        RECT 20.970 8.750 21.140 10.380 ;
        RECT 20.090 8.580 21.140 8.750 ;
        RECT 18.110 8.430 18.360 8.490 ;
        RECT 17.640 8.130 18.360 8.430 ;
        RECT 17.640 7.600 17.810 8.130 ;
        RECT 18.140 7.510 18.310 7.840 ;
        RECT 18.620 7.610 18.790 8.490 ;
        RECT 19.730 7.610 19.900 8.500 ;
        RECT 21.820 7.990 21.990 10.730 ;
        RECT 22.400 8.500 22.570 10.920 ;
        RECT 22.840 10.140 23.010 10.730 ;
        RECT 23.400 10.310 23.570 10.980 ;
        RECT 23.840 10.140 24.010 10.730 ;
        RECT 24.400 10.310 24.570 10.980 ;
        RECT 24.840 10.140 25.010 10.730 ;
        RECT 25.400 10.310 25.570 10.980 ;
        RECT 25.840 10.140 26.010 10.730 ;
        RECT 26.400 10.310 26.570 10.980 ;
        RECT 26.840 10.140 27.010 10.730 ;
        RECT 27.400 10.310 27.570 10.980 ;
        RECT 27.840 10.140 28.010 10.730 ;
        RECT 28.400 10.310 28.570 10.980 ;
        RECT 28.840 10.140 29.010 10.730 ;
        RECT 22.840 9.820 29.010 10.140 ;
        RECT 22.840 9.430 23.990 9.820 ;
        RECT 25.420 9.460 26.010 9.820 ;
        RECT 22.840 8.500 23.010 9.430 ;
        RECT 25.150 9.290 26.230 9.460 ;
        RECT 26.790 9.270 27.440 9.560 ;
        RECT 29.580 9.490 29.950 11.990 ;
        RECT 32.090 9.920 33.670 10.130 ;
        RECT 31.310 9.630 31.480 9.650 ;
        RECT 24.050 8.850 26.230 9.020 ;
        RECT 21.820 7.570 23.060 7.990 ;
        RECT 24.050 7.770 24.250 8.850 ;
        RECT 26.780 8.770 27.450 9.270 ;
        RECT 27.880 9.240 29.950 9.490 ;
        RECT 31.190 9.400 31.480 9.630 ;
        RECT 30.150 9.070 30.510 9.130 ;
        RECT 27.890 8.800 28.970 8.970 ;
        RECT 29.360 8.870 30.510 9.070 ;
        RECT 30.150 8.840 30.510 8.870 ;
        RECT 24.520 8.420 24.690 8.650 ;
        RECT 26.790 8.520 27.450 8.770 ;
        RECT 28.070 8.520 28.770 8.800 ;
        RECT 26.790 8.480 28.770 8.520 ;
        RECT 29.300 8.480 29.470 8.640 ;
        RECT 24.520 7.900 25.860 8.420 ;
        RECT 26.790 8.200 29.470 8.480 ;
        RECT 24.520 7.810 24.690 7.900 ;
        RECT 29.300 7.800 29.470 8.200 ;
        RECT 29.740 7.800 29.910 8.640 ;
        RECT 31.310 8.050 31.480 9.400 ;
        RECT 31.750 8.050 31.920 9.650 ;
        RECT 32.090 7.880 32.260 9.920 ;
        RECT 32.440 8.050 32.610 9.650 ;
        RECT 33.500 8.050 33.670 9.920 ;
        RECT 31.440 7.670 32.260 7.880 ;
        RECT 33.940 7.510 34.110 8.410 ;
        RECT 33.820 7.310 34.230 7.510 ;
        RECT 2.560 5.340 3.250 5.700 ;
        RECT 1.380 5.090 3.250 5.340 ;
        RECT 3.850 5.500 4.560 5.690 ;
        RECT 1.380 4.410 1.650 5.090 ;
        RECT 3.850 5.030 4.290 5.500 ;
        RECT 6.270 5.370 6.490 6.240 ;
        RECT 6.270 5.200 7.110 5.370 ;
        RECT 7.280 5.240 7.570 6.240 ;
        RECT 10.390 5.850 29.150 6.040 ;
        RECT 17.040 5.800 17.420 5.850 ;
        RECT 18.300 5.800 18.680 5.850 ;
        RECT 20.540 5.800 20.920 5.850 ;
        RECT 9.890 5.360 10.830 5.550 ;
        RECT 11.150 5.360 29.150 5.550 ;
        RECT 17.040 5.310 17.420 5.360 ;
        RECT 18.300 5.310 18.680 5.360 ;
        RECT 6.910 5.070 7.110 5.200 ;
        RECT 3.850 4.910 6.720 5.030 ;
        RECT 1.880 4.860 6.720 4.910 ;
        RECT 1.880 4.650 4.300 4.860 ;
        RECT 6.910 4.730 7.140 5.070 ;
        RECT 6.910 4.690 7.100 4.730 ;
        RECT 6.260 4.520 7.100 4.690 ;
        RECT 1.380 4.170 4.110 4.410 ;
        RECT 6.260 4.140 6.480 4.520 ;
        RECT 7.400 4.500 7.570 5.240 ;
        RECT 7.270 4.020 7.570 4.500 ;
        RECT 10.710 4.490 10.880 4.820 ;
        RECT 11.150 4.810 17.690 4.980 ;
        RECT 20.540 4.960 20.920 5.360 ;
        RECT 16.660 4.220 16.910 4.810 ;
        RECT 17.100 4.760 17.690 4.810 ;
        RECT 20.520 4.770 20.940 4.960 ;
        RECT 17.150 4.710 17.690 4.760 ;
        RECT 17.220 4.650 17.690 4.710 ;
        RECT 17.270 4.290 17.690 4.650 ;
        RECT 19.890 4.540 20.220 4.710 ;
        RECT 20.520 4.330 29.950 4.480 ;
        RECT 16.620 4.050 16.950 4.220 ;
        RECT 19.280 3.950 29.950 4.330 ;
        RECT 19.280 3.940 20.630 3.950 ;
        RECT 29.070 3.940 29.950 3.950 ;
        RECT 0.390 2.440 0.820 2.750 ;
        RECT 1.910 2.520 2.240 2.690 ;
        RECT 3.870 1.320 4.060 3.780 ;
        RECT 4.350 2.970 4.540 3.780 ;
        RECT 5.230 3.080 5.420 3.210 ;
        RECT 4.960 2.970 5.420 3.080 ;
        RECT 4.350 2.720 5.420 2.970 ;
        RECT 4.350 2.660 4.650 2.720 ;
        RECT 4.350 1.550 4.610 2.660 ;
        RECT 4.960 2.640 5.420 2.720 ;
        RECT 5.230 2.530 5.420 2.640 ;
        RECT 5.710 2.310 5.900 3.180 ;
        RECT 6.520 2.520 6.740 3.390 ;
        RECT 6.520 2.350 7.360 2.520 ;
        RECT 7.530 2.390 7.820 3.390 ;
        RECT 5.400 2.080 5.900 2.310 ;
        RECT 7.170 2.220 7.360 2.350 ;
        RECT 6.150 2.010 6.970 2.180 ;
        RECT 7.170 1.930 7.390 2.220 ;
        RECT 4.350 1.320 4.540 1.550 ;
        RECT 4.970 1.210 5.430 1.900 ;
        RECT 7.160 1.880 7.390 1.930 ;
        RECT 7.160 1.840 7.340 1.880 ;
        RECT 6.510 1.670 7.340 1.840 ;
        RECT 6.510 1.290 6.730 1.670 ;
        RECT 7.650 1.650 7.820 2.390 ;
        RECT 10.080 2.960 10.340 3.220 ;
        RECT 9.370 2.120 9.700 2.290 ;
        RECT 7.520 1.170 7.820 1.650 ;
        RECT 9.600 1.150 9.790 1.910 ;
        RECT 10.080 1.190 10.270 2.960 ;
        RECT 18.770 2.950 18.940 3.280 ;
        RECT 19.280 3.190 19.630 3.940 ;
        RECT 19.210 3.020 19.630 3.190 ;
        RECT 10.610 2.120 10.940 2.290 ;
        RECT 11.320 2.200 11.510 2.860 ;
        RECT 12.040 2.520 12.990 2.710 ;
        RECT 19.210 2.680 19.630 2.710 ;
        RECT 18.660 2.630 19.630 2.680 ;
        RECT 13.290 2.440 19.630 2.630 ;
        RECT 10.840 1.160 11.030 1.920 ;
        RECT 11.320 1.840 12.980 2.200 ;
        RECT 13.290 1.960 19.820 2.150 ;
        RECT 11.320 1.200 11.510 1.840 ;
        RECT 18.840 1.560 19.090 1.960 ;
        RECT 19.270 1.920 19.820 1.960 ;
        RECT 19.340 1.880 19.820 1.920 ;
        RECT 19.390 1.830 19.820 1.880 ;
        RECT 19.400 1.630 19.820 1.830 ;
        RECT 18.800 1.390 19.130 1.560 ;
        RECT 19.400 1.150 19.820 1.360 ;
      LAYER mcon ;
        RECT 9.320 11.400 9.490 11.570 ;
        RECT 10.400 11.480 10.570 11.650 ;
        RECT 11.060 11.380 11.230 11.550 ;
        RECT 12.040 10.830 12.210 11.000 ;
        RECT 13.330 10.770 13.500 10.940 ;
        RECT 16.060 12.350 16.230 12.530 ;
        RECT 16.980 11.370 17.150 11.540 ;
        RECT 17.590 11.380 17.760 11.550 ;
        RECT 21.820 11.590 21.990 11.760 ;
        RECT 22.070 10.980 22.240 11.150 ;
        RECT 29.170 10.980 29.340 11.150 ;
        RECT 19.480 10.640 19.650 10.810 ;
        RECT 3.710 9.120 3.880 9.290 ;
        RECT 2.070 8.470 2.240 8.640 ;
        RECT 2.730 8.570 2.900 8.740 ;
        RECT 3.680 7.650 3.850 7.820 ;
        RECT 5.000 9.180 5.170 9.350 ;
        RECT 7.720 9.140 7.890 9.310 ;
        RECT 8.650 8.580 8.820 8.750 ;
        RECT 9.260 8.570 9.430 8.740 ;
        RECT 9.760 8.580 9.930 8.750 ;
        RECT 7.730 7.590 7.900 7.770 ;
        RECT 14.120 9.120 14.290 9.290 ;
        RECT 12.480 8.470 12.650 8.640 ;
        RECT 13.140 8.570 13.310 8.740 ;
        RECT 14.090 7.650 14.260 7.820 ;
        RECT 15.410 9.180 15.580 9.350 ;
        RECT 18.130 9.140 18.300 9.310 ;
        RECT 19.060 8.580 19.230 8.750 ;
        RECT 19.670 8.570 19.840 8.740 ;
        RECT 20.170 8.580 20.340 8.750 ;
        RECT 18.140 7.590 18.310 7.770 ;
        RECT 27.040 9.310 27.210 9.480 ;
        RECT 31.220 9.430 31.390 9.600 ;
        RECT 27.040 8.840 27.210 9.010 ;
        RECT 30.190 8.860 30.480 9.110 ;
        RECT 22.880 7.700 23.050 7.870 ;
        RECT 24.080 7.970 24.250 8.140 ;
        RECT 25.580 7.960 25.800 8.160 ;
        RECT 29.740 8.030 29.910 8.200 ;
        RECT 31.750 9.430 31.920 9.600 ;
        RECT 32.440 8.590 32.610 8.760 ;
        RECT 21.480 5.860 21.650 6.030 ;
        RECT 21.820 5.860 21.990 6.030 ;
        RECT 10.710 4.570 10.880 4.740 ;
        RECT 19.970 4.540 20.140 4.710 ;
        RECT 29.580 4.170 29.750 4.340 ;
        RECT 0.450 2.480 0.760 2.700 ;
        RECT 1.990 2.520 2.160 2.690 ;
        RECT 3.880 1.700 4.050 1.870 ;
        RECT 4.440 2.690 4.610 2.860 ;
        RECT 6.210 2.010 6.380 2.180 ;
        RECT 5.100 1.460 5.270 1.630 ;
        RECT 10.130 3.000 10.300 3.170 ;
        RECT 18.770 3.030 18.940 3.200 ;
        RECT 9.450 2.120 9.620 2.290 ;
        RECT 9.610 1.570 9.780 1.740 ;
        RECT 9.610 1.230 9.780 1.400 ;
        RECT 10.690 2.120 10.860 2.290 ;
        RECT 10.850 1.580 11.020 1.750 ;
        RECT 10.850 1.240 11.020 1.410 ;
        RECT 19.530 1.180 19.700 1.350 ;
      LAYER met1 ;
        RECT 15.980 12.280 16.300 12.600 ;
        RECT 9.230 11.320 9.580 11.660 ;
        RECT 10.320 11.430 10.630 11.710 ;
        RECT 10.330 11.060 10.600 11.430 ;
        RECT 10.980 11.320 17.210 11.600 ;
        RECT 17.490 11.300 17.840 11.650 ;
        RECT 21.250 11.530 22.050 11.820 ;
        RECT 10.330 10.790 12.270 11.060 ;
        RECT 11.950 10.770 12.270 10.790 ;
        RECT 11.950 10.760 12.260 10.770 ;
        RECT 13.260 10.690 13.590 11.020 ;
        RECT 19.400 10.570 19.720 10.890 ;
        RECT 21.250 10.290 21.450 11.530 ;
        RECT 22.040 11.200 29.400 11.210 ;
        RECT 22.030 10.920 29.400 11.200 ;
        RECT 21.140 9.810 30.110 10.290 ;
        RECT 3.620 9.350 3.930 9.360 ;
        RECT 3.620 9.330 3.940 9.350 ;
        RECT 2.000 9.060 3.940 9.330 ;
        RECT 4.930 9.100 5.260 9.430 ;
        RECT 7.630 9.080 9.980 9.370 ;
        RECT 14.030 9.350 14.340 9.360 ;
        RECT 14.030 9.330 14.350 9.350 ;
        RECT 2.000 8.690 2.270 9.060 ;
        RECT 1.990 8.410 2.300 8.690 ;
        RECT 2.650 8.520 8.880 8.800 ;
        RECT 9.160 8.470 9.510 8.820 ;
        RECT 9.700 8.790 9.980 9.080 ;
        RECT 12.410 9.060 14.350 9.330 ;
        RECT 15.340 9.100 15.670 9.430 ;
        RECT 18.040 9.080 20.390 9.370 ;
        RECT 3.620 7.990 9.020 8.240 ;
        RECT 3.620 7.570 3.910 7.990 ;
        RECT 8.770 7.880 9.020 7.990 ;
        RECT 9.700 7.880 9.990 8.790 ;
        RECT 12.410 8.690 12.680 9.060 ;
        RECT 12.400 8.410 12.710 8.690 ;
        RECT 13.060 8.520 19.290 8.800 ;
        RECT 19.570 8.470 19.920 8.820 ;
        RECT 20.110 8.790 20.390 9.080 ;
        RECT 3.620 7.560 3.900 7.570 ;
        RECT 7.650 7.520 7.970 7.840 ;
        RECT 8.770 7.560 9.990 7.880 ;
        RECT 14.030 7.990 19.430 8.240 ;
        RECT 14.030 7.570 14.320 7.990 ;
        RECT 19.180 7.880 19.430 7.990 ;
        RECT 20.110 7.880 20.400 8.790 ;
        RECT 26.780 8.770 27.450 9.810 ;
        RECT 30.630 9.370 31.450 9.660 ;
        RECT 31.690 9.370 35.020 9.660 ;
        RECT 30.630 9.190 30.900 9.370 ;
        RECT 30.050 8.820 30.900 9.190 ;
        RECT 30.050 8.770 32.670 8.820 ;
        RECT 26.790 8.760 27.440 8.770 ;
        RECT 30.610 8.530 32.670 8.770 ;
        RECT 22.810 7.920 24.310 8.190 ;
        RECT 14.030 7.560 14.310 7.570 ;
        RECT 18.060 7.520 18.380 7.840 ;
        RECT 19.180 7.560 20.400 7.880 ;
        RECT 22.820 7.640 23.110 7.920 ;
        RECT 25.520 7.900 29.970 8.260 ;
        RECT 21.420 5.800 22.100 6.090 ;
        RECT 10.630 4.490 10.950 4.810 ;
        RECT 19.890 4.480 20.210 4.780 ;
        RECT 29.510 4.100 29.830 4.420 ;
        RECT 0.390 2.470 2.220 2.750 ;
        RECT 4.350 2.600 4.700 2.950 ;
        RECT 10.050 2.920 10.370 3.240 ;
        RECT 18.690 2.950 19.010 3.270 ;
        RECT 0.390 2.440 0.820 2.470 ;
        RECT 6.140 1.930 6.460 2.250 ;
        RECT 9.380 2.040 9.700 2.360 ;
        RECT 10.610 2.040 10.930 2.360 ;
        RECT 21.350 2.000 22.140 2.750 ;
        RECT 3.820 1.690 4.800 1.930 ;
        RECT 3.820 1.640 5.330 1.690 ;
        RECT 4.570 1.400 5.330 1.640 ;
        RECT 9.570 1.450 9.820 1.800 ;
        RECT 10.810 1.450 11.060 1.810 ;
        RECT 21.350 1.450 21.830 2.000 ;
        RECT 9.570 1.150 21.830 1.450 ;
      LAYER via ;
        RECT 16.010 12.310 16.270 12.570 ;
        RECT 9.260 11.350 9.540 11.630 ;
        RECT 17.530 11.350 17.790 11.610 ;
        RECT 13.290 10.720 13.560 10.990 ;
        RECT 19.430 10.600 19.690 10.860 ;
        RECT 4.960 9.130 5.230 9.400 ;
        RECT 9.200 8.510 9.460 8.770 ;
        RECT 15.370 9.130 15.640 9.400 ;
        RECT 19.610 8.510 19.870 8.770 ;
        RECT 7.680 7.550 7.940 7.810 ;
        RECT 34.730 9.390 34.990 9.650 ;
        RECT 18.090 7.550 18.350 7.810 ;
        RECT 21.600 5.800 21.860 6.060 ;
        RECT 10.660 4.520 10.920 4.780 ;
        RECT 19.920 4.490 20.180 4.750 ;
        RECT 29.540 4.130 29.800 4.390 ;
        RECT 10.080 2.950 10.340 3.210 ;
        RECT 18.720 2.980 18.980 3.240 ;
        RECT 4.380 2.630 4.670 2.920 ;
        RECT 6.170 1.960 6.430 2.220 ;
        RECT 9.410 2.070 9.670 2.330 ;
        RECT 10.640 2.070 10.900 2.330 ;
        RECT 21.480 2.200 22.020 2.560 ;
      LAYER met2 ;
        RECT 9.210 11.290 9.600 11.680 ;
        RECT 15.980 11.630 16.300 12.570 ;
        RECT 17.490 11.650 17.820 11.720 ;
        RECT 17.490 11.630 17.840 11.650 ;
        RECT 13.270 11.340 17.840 11.630 ;
        RECT 13.270 10.990 13.600 11.340 ;
        RECT 17.490 11.300 17.840 11.340 ;
        RECT 13.260 10.930 13.600 10.990 ;
        RECT 13.260 10.690 13.590 10.930 ;
        RECT 19.370 10.540 19.750 10.920 ;
        RECT 4.930 9.190 5.260 9.430 ;
        RECT 15.340 9.190 15.670 9.430 ;
        RECT 4.930 9.130 5.270 9.190 ;
        RECT 15.340 9.130 15.680 9.190 ;
        RECT 4.940 8.780 5.270 9.130 ;
        RECT 9.160 8.780 9.510 8.820 ;
        RECT 4.940 8.490 9.510 8.780 ;
        RECT 15.350 8.780 15.680 9.130 ;
        RECT 19.570 8.780 19.920 8.820 ;
        RECT 15.350 8.490 19.920 8.780 ;
        RECT 7.650 7.550 7.970 8.490 ;
        RECT 9.160 8.470 9.510 8.490 ;
        RECT 9.160 8.400 9.490 8.470 ;
        RECT 18.060 7.550 18.380 8.490 ;
        RECT 19.570 8.470 19.920 8.490 ;
        RECT 19.570 8.400 19.900 8.470 ;
        RECT 34.700 6.860 35.020 9.660 ;
        RECT 30.320 6.540 35.020 6.860 ;
        RECT 10.510 4.790 10.950 4.810 ;
        RECT 9.270 4.490 10.950 4.790 ;
        RECT 9.270 4.430 10.940 4.490 ;
        RECT 17.370 4.460 20.210 4.780 ;
        RECT 9.270 3.180 9.590 4.430 ;
        RECT 17.370 3.460 17.840 4.460 ;
        RECT 4.350 2.920 4.700 2.950 ;
        RECT 4.350 2.650 6.410 2.920 ;
        RECT 8.680 2.870 9.590 3.180 ;
        RECT 10.050 3.060 17.840 3.460 ;
        RECT 10.050 2.920 10.370 3.060 ;
        RECT 18.140 2.950 19.010 3.270 ;
        RECT 4.350 2.600 4.700 2.650 ;
        RECT 6.150 2.250 6.410 2.650 ;
        RECT 9.270 2.360 9.590 2.870 ;
        RECT 6.140 1.930 6.460 2.250 ;
        RECT 9.270 2.040 9.700 2.360 ;
        RECT 10.430 2.070 10.930 2.360 ;
        RECT 10.430 1.560 10.760 2.070 ;
        RECT 18.140 1.560 18.510 2.950 ;
        RECT 21.450 2.170 22.060 6.090 ;
        RECT 30.320 4.420 30.670 6.540 ;
        RECT 29.510 4.100 30.670 4.420 ;
        RECT 10.430 1.550 18.510 1.560 ;
        RECT 8.680 1.190 18.510 1.550 ;
      LAYER via2 ;
        RECT 9.260 11.340 9.540 11.620 ;
        RECT 19.420 10.590 19.700 10.870 ;
      LAYER met3 ;
        RECT 8.910 11.290 9.600 11.680 ;
        RECT 8.910 10.610 9.260 11.290 ;
        RECT 19.370 10.850 19.750 10.920 ;
        RECT 19.370 10.610 19.790 10.850 ;
        RECT 8.910 10.260 19.790 10.610 ;
  END
END avsdpll
END LIBRARY
