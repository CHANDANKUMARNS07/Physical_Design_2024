VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO avsddac
  CLASS BLOCK ;
  FOREIGN avsddac ;
  ORIGIN -136.770 -613.050 ;
  SIZE 1193.570 BY 562.310 ;
  PIN D[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1150.220 613.050 1151.250 755.620 ;
    END
  END D[9]
  PIN D[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1117.200 613.050 1117.850 709.180 ;
    END
  END D[8]
  PIN D[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1096.950 613.050 1097.260 619.510 ;
    END
  END D[7]
  PIN D[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1078.220 613.050 1079.660 614.760 ;
    END
  END D[6]
  PIN D[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 226.250 1174.740 228.070 1175.360 ;
    END
  END D[5]
  PIN D[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 209.700 1174.310 211.150 1175.360 ;
    END
  END D[4]
  PIN D[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met1 ;
        RECT 432.010 1168.710 433.190 1175.360 ;
    END
  END D[3]
  PIN D[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 178.380 1174.680 180.110 1175.360 ;
    END
  END D[2]
  PIN D[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 160.760 1172.150 162.090 1175.360 ;
    END
  END D[1]
  PIN D[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 145.960 1172.220 146.570 1175.360 ;
    END
  END D[0]
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 152.670 1171.410 154.120 1175.360 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met2 ;
        RECT 136.770 873.200 144.500 873.520 ;
    END
  END VGND
  PIN VREFH
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 142.900 1170.680 143.170 1175.360 ;
    END
  END VREFH
  PIN OUT
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met4 ;
        RECT 1172.680 1127.710 1173.730 1175.360 ;
    END
  END OUT
  OBS
      LAYER li1 ;
        RECT 136.770 1170.510 142.730 1175.360 ;
        RECT 143.340 1172.050 145.790 1175.360 ;
        RECT 146.740 1172.050 160.590 1175.360 ;
        RECT 143.340 1171.980 160.590 1172.050 ;
        RECT 162.260 1174.510 178.210 1175.360 ;
        RECT 180.280 1174.510 209.530 1175.360 ;
        RECT 162.260 1174.140 209.530 1174.510 ;
        RECT 211.320 1174.570 226.080 1175.360 ;
        RECT 228.240 1174.570 1164.190 1175.360 ;
        RECT 211.320 1174.140 1164.190 1174.570 ;
        RECT 162.260 1171.980 1164.190 1174.140 ;
        RECT 143.340 1170.510 1164.190 1171.980 ;
        RECT 136.770 755.790 1164.190 1170.510 ;
        RECT 136.770 709.350 1150.050 755.790 ;
        RECT 136.770 619.680 1117.030 709.350 ;
        RECT 136.770 614.930 1096.780 619.680 ;
        RECT 136.770 613.050 1078.050 614.930 ;
        RECT 1079.830 613.050 1096.780 614.930 ;
        RECT 1097.430 613.050 1117.030 619.680 ;
        RECT 1118.020 613.050 1150.050 709.350 ;
        RECT 1151.420 613.050 1164.190 755.790 ;
      LAYER met1 ;
        RECT 140.750 1168.430 431.730 1175.360 ;
        RECT 433.470 1168.430 1313.360 1175.360 ;
        RECT 140.750 613.050 1313.360 1168.430 ;
      LAYER met2 ;
        RECT 143.250 873.800 1165.380 1172.180 ;
        RECT 144.780 872.920 1165.380 873.800 ;
        RECT 143.250 641.910 1165.380 872.920 ;
      LAYER met3 ;
        RECT 146.990 647.680 1330.340 1169.670 ;
      LAYER met4 ;
        RECT 147.000 1171.010 152.270 1175.050 ;
        RECT 154.520 1171.010 1172.280 1175.050 ;
        RECT 147.000 1127.310 1172.280 1171.010 ;
        RECT 1174.130 1127.310 1188.200 1175.050 ;
        RECT 147.000 648.540 1188.200 1127.310 ;
  END
END avsddac
END LIBRARY
